`define IOB_IBEX_AXI_ID_W 0
`define IOB_IBEX_AXI_ADDR_W 32
`define IOB_IBEX_AXI_DATA_W 32
`define IOB_IBEX_AXI_LEN_W 8
`define IOB_IBEX_IBEX_ADDR_W 32
`define IOB_IBEX_IBEX_DATA_W 32
`define IOB_IBEX_IBEX_INTG_DATA_W 7
