`ifndef FATORI_SELFTEST_SVH
`define FATORI_SELFTEST_SVH


`endif // FATORI_SELFTEST_SVH