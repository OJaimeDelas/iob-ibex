`ifndef FATORI_PBLOCKS_SVH
`define FATORI_PBLOCKS_SVH

`define KEEP_ALU (* keep_hierarchy = "true" *)
`define KEEP_MULTIPLIER (* keep_hierarchy = "true" *)
`define KEEP_CONTROLLER (* keep_hierarchy = "true" *)
`define KEEP_DECODER (* keep_hierarchy = "true" *)
`define KEEP_LSU (* keep_hierarchy = "true" *)
`define KEEP_IF_STAGE (* keep_hierarchy = "true" *)
`define KEEP_ID_STAGE (* keep_hierarchy = "true" *)
`define KEEP_WB_STAGE (* keep_hierarchy = "true" *)
`define KEEP_PREFETCH_BUFFER (* keep_hierarchy = "true" *)
`define KEEP_BRANCH_PREDICT (* keep_hierarchy = "true" *)
`define KEEP_FAULT_MGR (* keep_hierarchy = "true" *)

`endif // FATORI_PBLOCKS_SVH